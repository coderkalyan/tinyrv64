module dut_harness ();
    register_file rf;
    decoder id;
    alu alu;
endmodule
